`timescale 1ns / 1ps
/*
To test the Entire Decode Stage 
*/
module Decode_Stage_tb();
    
endmodule