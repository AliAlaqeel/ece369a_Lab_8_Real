`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369 - Computer Architecture
// 
// Module - ALU32Bit.v
// Description - 32-Bit wide arithmetic logic unit (ALU).
//
// INPUTS:-
// ALUControl: N-Bit input control bits to select an ALU operation.
// A: 32-Bit input port A.
// B: 32-Bit input port B.
//
// OUTPUTS:-
// ALUResult: 32-Bit ALU result output.
// ZERO: 1-Bit output flag. 
//
// FUNCTIONALITY:-
// Design a 32-Bit ALU, so that it supports all arithmetic operations 
// needed by the MIPS instructions given in Labs5-8.docx document. 
//   The 'ALUResult' will output the corresponding result of the operation 
//   based on the 32-Bit inputs, 'A', and 'B'. 
//   The 'Zero' flag is high when 'ALUResult' is '0'. 
//   The 'ALUControl' signal should determine the function of the ALU 
//   You need to determine the bitwidth of the ALUControl signal based on the number of 
//   operations needed to support. 
////////////////////////////////////////////////////////////////////////////////

module ALU32Bit(ALUControl, A, B, ALUResult, Zero);

	input [3:0] ALUControl; // control bits for ALU operation
                                // you need to adjust the bitwidth as needed
	input signed [31:0] A, B;	    // inputs

	output reg [31:0] ALUResult;	// answer
	output reg Zero;	    // Zero=1 if ALUResult == 0

    /* Please fill in the implementation here... */
	always@(*)begin
		case(ALUControl)
			0: ALUResult <= A + B;	//Add, Addi, Loads & Stores
			1: ALUResult <= A - B;	//Sub
			2: ALUResult <= A * B;	//Mul
			3: ALUResult <= A & B;	//And
			4: ALUResult <= A | B;	//Or
			5: ALUResult <= ~(A | B);	//NOr
			6: ALUResult <= A <<< $unsigned(B);	//Shift left
			7: ALUResult <= A >>> $unsigned(B);	//Shift right
			8: ALUResult <= A ^ B;	//Xor
			9: begin				//Slt, Slti
				if(A < B) ALUResult <= 1;
				else ALUResult <= 0;
			end
			10: ALUResult <= 0;		//Jumps
			11: ALUResult <= A;		//Pass Value of A
			default: ALUResult <= 32'd2147483647;
		endcase
	end

	always@(*)begin
		if(ALUResult == 0) Zero <= 1;
		else Zero <= 0;
	end
endmodule
